module(
    input [8:0] IN,
    output [24:0] OUT
);

always@(*) begin
    case(IN):
        3: OUT = 9686330;
        4: OUT = 8388608;
        5: OUT = 7502999;
        6: OUT = 6849269;
        7: OUT = 6341191;
        8: OUT = 5931641;
        9: OUT = 5592405;
        10: OUT = 5305421;
        11: OUT = 5058520;
        12: OUT = 4843165;
        13: OUT = 4653162;
        14: OUT = 4483899;
        15: OUT = 4331858;
        16: OUT = 4194304;
        17: OUT = 4069072;
        18: OUT = 3954427;
        19: OUT = 3848957;
        20: OUT = 3751499;
        21: OUT = 3661088;
        22: OUT = 3576914;
        23: OUT = 3498291;
        24: OUT = 3424634;
        25: OUT = 3355443;
        26: OUT = 3290282;
        27: OUT = 3228776;
        28: OUT = 3170595;
        29: OUT = 3115450;
        30: OUT = 3063086;
        31: OUT = 3013276;
        32: OUT = 2965820;
        33: OUT = 2920538;
        34: OUT = 2877268;
        35: OUT = 2835867;
        36: OUT = 2796202;
        37: OUT = 2758157;
        38: OUT = 2721623;
        39: OUT = 2686504;
        40: OUT = 2652710;
        41: OUT = 2620160;
        42: OUT = 2588780;
        43: OUT = 2558501;
        44: OUT = 2529260;
        45: OUT = 2500999;
        46: OUT = 2473665;
        47: OUT = 2447208;
        48: OUT = 2421582;
        49: OUT = 2396745;
        50: OUT = 2372656;
        51: OUT = 2349280;
        52: OUT = 2326581;
        53: OUT = 2304527;
        54: OUT = 2283089;
        55: OUT = 2262239;
        56: OUT = 2241949;
        57: OUT = 2222196;
        58: OUT = 2202956;
        59: OUT = 2184207;
        60: OUT = 2165929;
        61: OUT = 2148102;
        62: OUT = 2130708;
        63: OUT = 2113730;
        64: OUT = 2097152;
        65: OUT = 2080957;
        66: OUT = 2065132;
        67: OUT = 2049663;
        68: OUT = 2034536;
        69: OUT = 2019739;
        70: OUT = 2005260;
        71: OUT = 1991089;
        72: OUT = 1977213;
        73: OUT = 1963624;
        74: OUT = 1950311;
        75: OUT = 1937266;
        76: OUT = 1924478;
        77: OUT = 1911941;
        78: OUT = 1899645;
        79: OUT = 1887584;
        80: OUT = 1875749;
        81: OUT = 1864135;
        82: OUT = 1852733;
        83: OUT = 1841538;
        84: OUT = 1830544;
        85: OUT = 1819744;
        86: OUT = 1809133;
        87: OUT = 1798706;
        88: OUT = 1788457;
        89: OUT = 1778381;
        90: OUT = 1768473;
        91: OUT = 1758730;
        92: OUT = 1749145;
        93: OUT = 1739716;
        94: OUT = 1730437;
        95: OUT = 1721306;
        96: OUT = 1712317;
        97: OUT = 1703468;
        98: OUT = 1694754;
        99: OUT = 1686173;
        100: OUT = 1677721;
        101: OUT = 1669395;
        102: OUT = 1661191;
        103: OUT = 1653108;
        104: OUT = 1645141;
        105: OUT = 1637288;
        106: OUT = 1629547;
        107: OUT = 1621914;
        108: OUT = 1614388;
        109: OUT = 1606965;
        110: OUT = 1599644;
        111: OUT = 1592422;
        112: OUT = 1585297;
        113: OUT = 1578267;
        114: OUT = 1571330;
        115: OUT = 1564483;
        116: OUT = 1557725;
        117: OUT = 1551054;
        118: OUT = 1544467;
        119: OUT = 1537964;
        120: OUT = 1531543;
        121: OUT = 1525201;
        122: OUT = 1518937;
        123: OUT = 1512750;
        124: OUT = 1506638;
        125: OUT = 1500599;
        126: OUT = 1494633;
        127: OUT = 1488737;
        128: OUT = 1482910;
        129: OUT = 1477151;
        130: OUT = 1471459;
        131: OUT = 1465832;
        132: OUT = 1460269;
        133: OUT = 1454769;
        134: OUT = 1449330;
        135: OUT = 1443952;
        136: OUT = 1438634;
        137: OUT = 1433374;
        138: OUT = 1428171;
        139: OUT = 1423024;
        140: OUT = 1417933;
        141: OUT = 1412896;
        142: OUT = 1407912;
        143: OUT = 1402981;
        144: OUT = 1398101;
        145: OUT = 1393271;
        146: OUT = 1388492;
        147: OUT = 1383761;
        148: OUT = 1379078;
        149: OUT = 1374443;
        150: OUT = 1369853;
        151: OUT = 1365310;
        152: OUT = 1360811;
        153: OUT = 1356357;
        154: OUT = 1351946;
        155: OUT = 1347578;
        156: OUT = 1343252;
        157: OUT = 1338967;
        158: OUT = 1334723;
        159: OUT = 1330519;
        160: OUT = 1326355;
        161: OUT = 1322229;
        162: OUT = 1318142;
        163: OUT = 1314092;
        164: OUT = 1310080;
        165: OUT = 1306104;
        166: OUT = 1302164;
        167: OUT = 1298259;
        168: OUT = 1294390;
        169: OUT = 1290555;
        170: OUT = 1286753;
        171: OUT = 1282985;
        172: OUT = 1279250;
        173: OUT = 1275548;
        174: OUT = 1271877;
        175: OUT = 1268238;
        176: OUT = 1264630;
        177: OUT = 1261052;
        178: OUT = 1257505;
        179: OUT = 1253987;
        180: OUT = 1250499;
        181: OUT = 1247040;
        182: OUT = 1243609;
        183: OUT = 1240207;
        184: OUT = 1236832;
        185: OUT = 1233485;
        186: OUT = 1230165;
        187: OUT = 1226871;
        188: OUT = 1223604;
        189: OUT = 1220362;
        190: OUT = 1217147;
        191: OUT = 1213956;
        192: OUT = 1210791;
        193: OUT = 1207650;
        194: OUT = 1204533;
        195: OUT = 1201441;
        196: OUT = 1198372;
        197: OUT = 1195327;
        198: OUT = 1192304;
        199: OUT = 1189305;
        200: OUT = 1186328;
        201: OUT = 1183373;
        202: OUT = 1180440;
        203: OUT = 1177529;
        204: OUT = 1174640;
        205: OUT = 1171771;
        206: OUT = 1168924;
        207: OUT = 1166097;
        208: OUT = 1163290;
        209: OUT = 1160504;
        210: OUT = 1157737;
        211: OUT = 1154991;
        212: OUT = 1152263;
        213: OUT = 1149555;
        214: OUT = 1146866;
        215: OUT = 1144196;
        216: OUT = 1141544;
        217: OUT = 1138911;
        218: OUT = 1136296;
        219: OUT = 1133699;
        220: OUT = 1131119;
        221: OUT = 1128557;
        222: OUT = 1126013;
        223: OUT = 1123485;
        224: OUT = 1120974;
        225: OUT = 1118481;
        226: OUT = 1116003;
        227: OUT = 1113542;
        228: OUT = 1111098;
        229: OUT = 1108669;
        230: OUT = 1106256;
        231: OUT = 1103859;
        232: OUT = 1101478;
        233: OUT = 1099111;
        234: OUT = 1096760;
        235: OUT = 1094424;
        236: OUT = 1092103;
        237: OUT = 1089797;
        238: OUT = 1087505;
        239: OUT = 1085227;
        240: OUT = 1082964;
        241: OUT = 1080715;
        242: OUT = 1078480;
        243: OUT = 1076258;
        244: OUT = 1074051;
        245: OUT = 1071857;
        246: OUT = 1069676;
        247: OUT = 1067508;
        248: OUT = 1065354;
        249: OUT = 1063212;
        250: OUT = 1061084;
        251: OUT = 1058968;
        252: OUT = 1056865;
        253: OUT = 1054774;
        254: OUT = 1052696;
        255: OUT = 1050630;
        256: OUT = 1048576;
        257: OUT = 1046533;
        258: OUT = 1044503;
        259: OUT = 1042485;
        260: OUT = 1040478;
        261: OUT = 1038483;
        262: OUT = 1036499;
        263: OUT = 1034527;
        264: OUT = 1032566;
        265: OUT = 1030616;
        266: OUT = 1028677;
        267: OUT = 1026748;
        268: OUT = 1024831;
        269: OUT = 1022924;
        270: OUT = 1021028;
        271: OUT = 1019143;
        272: OUT = 1017268;
        273: OUT = 1015403;
        274: OUT = 1013548;
        275: OUT = 1011704;
        276: OUT = 1009869;
        277: OUT = 1008045;
        278: OUT = 1006230;
        279: OUT = 1004425;
        280: OUT = 1002630;
        281: OUT = 1000844;
        282: OUT = 999068;
        283: OUT = 997301;
        284: OUT = 995544;
        285: OUT = 993796;
        286: OUT = 992057;
        287: OUT = 990327;
        288: OUT = 988606;
        289: OUT = 986895;
        290: OUT = 985192;
        291: OUT = 983497;
        292: OUT = 981812;
        293: OUT = 980135;
        294: OUT = 978467;
        295: OUT = 976807;
        296: OUT = 975155;
        297: OUT = 973512;
        298: OUT = 971878;
        299: OUT = 970251;
        300: OUT = 968633;
        301: OUT = 967022;
        302: OUT = 965420;
        303: OUT = 963825;
        304: OUT = 962239;
        305: OUT = 960660;
        306: OUT = 959089;
        307: OUT = 957526;
        308: OUT = 955970;
        309: OUT = 954422;
        310: OUT = 952881;
        311: OUT = 951348;
        312: OUT = 949822;
        313: OUT = 948304;
        314: OUT = 946793;
        315: OUT = 945289;
        316: OUT = 943792;
        317: OUT = 942302;
        318: OUT = 940819;
        319: OUT = 939343;
        320: OUT = 937874;
        321: OUT = 936412;
        322: OUT = 934957;
        323: OUT = 933509;
        324: OUT = 932067;
        325: OUT = 930632;
        326: OUT = 929204;
        327: OUT = 927782;
        328: OUT = 926366;
        329: OUT = 924957;
        330: OUT = 923555;
        331: OUT = 922159;
        332: OUT = 920769;
        333: OUT = 919385;
        334: OUT = 918008;
        335: OUT = 916637;
        336: OUT = 915272;
        337: OUT = 913913;
        338: OUT = 912560;
        339: OUT = 911213;
        340: OUT = 909872;
        341: OUT = 908537;
        342: OUT = 907207;
        343: OUT = 905884;
        344: OUT = 904566;
        345: OUT = 903254;
        346: OUT = 901948;
        347: OUT = 900648;
        348: OUT = 899353;
        349: OUT = 898063;
        350: OUT = 896779;
        351: OUT = 895501;
        352: OUT = 894228;
        353: OUT = 892961;
        354: OUT = 891698;
        355: OUT = 890442;
        356: OUT = 889190;
        357: OUT = 887944;
        358: OUT = 886703;
        359: OUT = 885467;
        360: OUT = 884236;
        361: OUT = 883011;
        362: OUT = 881790;
        363: OUT = 880575;
        364: OUT = 879365;
        365: OUT = 878159;
        366: OUT = 876959;
        367: OUT = 875763;
        368: OUT = 874572;
        369: OUT = 873386;
        370: OUT = 872205;
        371: OUT = 871029;
        372: OUT = 869858;
        373: OUT = 868691;
        374: OUT = 867529;
        375: OUT = 866371;
        376: OUT = 865218;
        377: OUT = 864070;
        378: OUT = 862926;
        379: OUT = 861787;
        380: OUT = 860653;
        381: OUT = 859522;
        382: OUT = 858397;
        383: OUT = 857275;
    endcase

end

endmodule