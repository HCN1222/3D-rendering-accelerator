
module controller(





);




endmodule