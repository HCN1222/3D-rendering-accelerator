


module vertice_shader(








);


    GetMVP GetMVP(
	
	
	
	);
	
	
	matrix_multiplication matrix_multiplication(
	
	
	
	);
	
	
	DO_NDC DO_NDC(
	
	
	
	
	);
	
	ChangeToScreen ChangeToScreen(
	
	
	
	);


endmodule


