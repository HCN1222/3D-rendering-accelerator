module NDC(
    input clk,
    input signed [23:0] x, //
    input signed [23:0] y,
    input signed [23:0] w,
    output signed reg [23:0] normalized_x,
    output signed reg [23:0] normalized_y,
);



endmodule