
module Rasterization(





);


    InTriangle InTriangle(
	
	
	
	
	);
	
	
	GetColorDepth GetColorDepth(
	
	
	
	
	
	);

endmodule
