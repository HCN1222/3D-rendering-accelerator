module dot_product(
    // input: 4Q20
    input [24:0] x1,
    input [24:0] y1,
    input [24:0] z1,

    input [24:0] x2,
    input [24:0] y2,
    input [24:0] z2,
    // output 
    output [24:0] out
);


endmodule